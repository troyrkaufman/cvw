 // specialCases.sv

 module specCase(input logic [15:0] x, y, z, product, sum,
                output logic [15:0] specAns
                output logic        of);
    // Is this just a string of if statements with a variety of inputs coming from the fmamult and fmaadd modules
   
   // 

    if () begin  end
    else if () begin  end
    else if () begin  end
    else if () begin  end
    else if () begin  end
    else if () begin  end
    else if () begin  end
    else        begin  end
 endmodule
